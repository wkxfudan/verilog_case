module not_gate(a,out);
       input wire a;
       output wire out;
       assign out=~a;

endmodule